`timescale 10ns / 1ps
module PRIORITY_ENCODER_4_2_tb();
reg [3:0] x;
wire [1:0] y;
PRIORITY_ENCODER_4_2 dut(.x(x), .y(y));
initial begin
x=4'b0000;#10
x=4'b0001;#10
x=4'b0010;#10
x=4'b0011;#10
x=4'b0100;#10
x=4'b0101;#10
x=4'b0110;#10
x=4'b0111;#10
x=4'b1000;#10
x=4'b1001;#10
x=4'b1010;#10
x=4'b1011;#10
x=4'b1100;#10
x=4'b1101;#10
x=4'b1110;#10
x=4'b1111;
end 
endmodule
